library verilog;
use verilog.vl_types.all;
entity tb_gfmul_v2 is
end tb_gfmul_v2;
