module gfmul(
//input [0:127] iR,
input [0:127] iCtext,
input [0:127] iHashkey,
output [0:127] oResult
);

// reg [0:127] Z;
// reg [0:127] V;
// integer idx;

// always @(*) begin
	// Z = 128'd0;
	// V = iHashkey;

	// for(idx = 0; idx <= 127; idx = idx + 1) begin
		// if(iCtext[idx])	Z = Z ^ V;
		// else			Z = Z;
		
		// if(~V[127])			V = {1'b0, V[0:126]}; // V = V >> 1;
		// else				V = {1'b0, V[0:126]} ^ {8'b11100001, 120'd0}; // V = V >> 1;
	// end
// end

// assign oResult = Z;


wire [0:127] Z [1:128];
wire [0:127] V [0:127];

wire [0:127] iR;
assign iR = {8'b1110_0001, 120'd0};

assign V[0] = iHashkey;
assign V[1] = {1'b0, V[0][0:126]} ^ (iR & {128{V[0][127]}});
assign V[2] = {1'b0, V[1][0:126]} ^ (iR & {128{V[1][127]}});
assign V[3] = {1'b0, V[2][0:126]} ^ (iR & {128{V[2][127]}});
assign V[4] = {1'b0, V[3][0:126]} ^ (iR & {128{V[3][127]}});
assign V[5] = {1'b0, V[4][0:126]} ^ (iR & {128{V[4][127]}});
assign V[6] = {1'b0, V[5][0:126]} ^ (iR & {128{V[5][127]}});
assign V[7] = {1'b0, V[6][0:126]} ^ (iR & {128{V[6][127]}});
assign V[8] = {1'b0, V[7][0:126]} ^ (iR & {128{V[7][127]}});
assign V[9] = {1'b0, V[8][0:126]} ^ (iR & {128{V[8][127]}});
assign V[10] = {1'b0, V[9][0:126]} ^ (iR & {128{V[9][127]}});
assign V[11] = {1'b0, V[10][0:126]} ^ (iR & {128{V[10][127]}});
assign V[12] = {1'b0, V[11][0:126]} ^ (iR & {128{V[11][127]}});
assign V[13] = {1'b0, V[12][0:126]} ^ (iR & {128{V[12][127]}});
assign V[14] = {1'b0, V[13][0:126]} ^ (iR & {128{V[13][127]}});
assign V[15] = {1'b0, V[14][0:126]} ^ (iR & {128{V[14][127]}});
assign V[16] = {1'b0, V[15][0:126]} ^ (iR & {128{V[15][127]}});
assign V[17] = {1'b0, V[16][0:126]} ^ (iR & {128{V[16][127]}});
assign V[18] = {1'b0, V[17][0:126]} ^ (iR & {128{V[17][127]}});
assign V[19] = {1'b0, V[18][0:126]} ^ (iR & {128{V[18][127]}});
assign V[20] = {1'b0, V[19][0:126]} ^ (iR & {128{V[19][127]}});
assign V[21] = {1'b0, V[20][0:126]} ^ (iR & {128{V[20][127]}});
assign V[22] = {1'b0, V[21][0:126]} ^ (iR & {128{V[21][127]}});
assign V[23] = {1'b0, V[22][0:126]} ^ (iR & {128{V[22][127]}});
assign V[24] = {1'b0, V[23][0:126]} ^ (iR & {128{V[23][127]}});
assign V[25] = {1'b0, V[24][0:126]} ^ (iR & {128{V[24][127]}});
assign V[26] = {1'b0, V[25][0:126]} ^ (iR & {128{V[25][127]}});
assign V[27] = {1'b0, V[26][0:126]} ^ (iR & {128{V[26][127]}});
assign V[28] = {1'b0, V[27][0:126]} ^ (iR & {128{V[27][127]}});
assign V[29] = {1'b0, V[28][0:126]} ^ (iR & {128{V[28][127]}});
assign V[30] = {1'b0, V[29][0:126]} ^ (iR & {128{V[29][127]}});
assign V[31] = {1'b0, V[30][0:126]} ^ (iR & {128{V[30][127]}});
assign V[32] = {1'b0, V[31][0:126]} ^ (iR & {128{V[31][127]}});
assign V[33] = {1'b0, V[32][0:126]} ^ (iR & {128{V[32][127]}});
assign V[34] = {1'b0, V[33][0:126]} ^ (iR & {128{V[33][127]}});
assign V[35] = {1'b0, V[34][0:126]} ^ (iR & {128{V[34][127]}});
assign V[36] = {1'b0, V[35][0:126]} ^ (iR & {128{V[35][127]}});
assign V[37] = {1'b0, V[36][0:126]} ^ (iR & {128{V[36][127]}});
assign V[38] = {1'b0, V[37][0:126]} ^ (iR & {128{V[37][127]}});
assign V[39] = {1'b0, V[38][0:126]} ^ (iR & {128{V[38][127]}});
assign V[40] = {1'b0, V[39][0:126]} ^ (iR & {128{V[39][127]}});
assign V[41] = {1'b0, V[40][0:126]} ^ (iR & {128{V[40][127]}});
assign V[42] = {1'b0, V[41][0:126]} ^ (iR & {128{V[41][127]}});
assign V[43] = {1'b0, V[42][0:126]} ^ (iR & {128{V[42][127]}});
assign V[44] = {1'b0, V[43][0:126]} ^ (iR & {128{V[43][127]}});
assign V[45] = {1'b0, V[44][0:126]} ^ (iR & {128{V[44][127]}});
assign V[46] = {1'b0, V[45][0:126]} ^ (iR & {128{V[45][127]}});
assign V[47] = {1'b0, V[46][0:126]} ^ (iR & {128{V[46][127]}});
assign V[48] = {1'b0, V[47][0:126]} ^ (iR & {128{V[47][127]}});
assign V[49] = {1'b0, V[48][0:126]} ^ (iR & {128{V[48][127]}});
assign V[50] = {1'b0, V[49][0:126]} ^ (iR & {128{V[49][127]}});
assign V[51] = {1'b0, V[50][0:126]} ^ (iR & {128{V[50][127]}});
assign V[52] = {1'b0, V[51][0:126]} ^ (iR & {128{V[51][127]}});
assign V[53] = {1'b0, V[52][0:126]} ^ (iR & {128{V[52][127]}});
assign V[54] = {1'b0, V[53][0:126]} ^ (iR & {128{V[53][127]}});
assign V[55] = {1'b0, V[54][0:126]} ^ (iR & {128{V[54][127]}});
assign V[56] = {1'b0, V[55][0:126]} ^ (iR & {128{V[55][127]}});
assign V[57] = {1'b0, V[56][0:126]} ^ (iR & {128{V[56][127]}});
assign V[58] = {1'b0, V[57][0:126]} ^ (iR & {128{V[57][127]}});
assign V[59] = {1'b0, V[58][0:126]} ^ (iR & {128{V[58][127]}});
assign V[60] = {1'b0, V[59][0:126]} ^ (iR & {128{V[59][127]}});
assign V[61] = {1'b0, V[60][0:126]} ^ (iR & {128{V[60][127]}});
assign V[62] = {1'b0, V[61][0:126]} ^ (iR & {128{V[61][127]}});
assign V[63] = {1'b0, V[62][0:126]} ^ (iR & {128{V[62][127]}});
assign V[64] = {1'b0, V[63][0:126]} ^ (iR & {128{V[63][127]}});
assign V[65] = {1'b0, V[64][0:126]} ^ (iR & {128{V[64][127]}});
assign V[66] = {1'b0, V[65][0:126]} ^ (iR & {128{V[65][127]}});
assign V[67] = {1'b0, V[66][0:126]} ^ (iR & {128{V[66][127]}});
assign V[68] = {1'b0, V[67][0:126]} ^ (iR & {128{V[67][127]}});
assign V[69] = {1'b0, V[68][0:126]} ^ (iR & {128{V[68][127]}});
assign V[70] = {1'b0, V[69][0:126]} ^ (iR & {128{V[69][127]}});
assign V[71] = {1'b0, V[70][0:126]} ^ (iR & {128{V[70][127]}});
assign V[72] = {1'b0, V[71][0:126]} ^ (iR & {128{V[71][127]}});
assign V[73] = {1'b0, V[72][0:126]} ^ (iR & {128{V[72][127]}});
assign V[74] = {1'b0, V[73][0:126]} ^ (iR & {128{V[73][127]}});
assign V[75] = {1'b0, V[74][0:126]} ^ (iR & {128{V[74][127]}});
assign V[76] = {1'b0, V[75][0:126]} ^ (iR & {128{V[75][127]}});
assign V[77] = {1'b0, V[76][0:126]} ^ (iR & {128{V[76][127]}});
assign V[78] = {1'b0, V[77][0:126]} ^ (iR & {128{V[77][127]}});
assign V[79] = {1'b0, V[78][0:126]} ^ (iR & {128{V[78][127]}});
assign V[80] = {1'b0, V[79][0:126]} ^ (iR & {128{V[79][127]}});
assign V[81] = {1'b0, V[80][0:126]} ^ (iR & {128{V[80][127]}});
assign V[82] = {1'b0, V[81][0:126]} ^ (iR & {128{V[81][127]}});
assign V[83] = {1'b0, V[82][0:126]} ^ (iR & {128{V[82][127]}});
assign V[84] = {1'b0, V[83][0:126]} ^ (iR & {128{V[83][127]}});
assign V[85] = {1'b0, V[84][0:126]} ^ (iR & {128{V[84][127]}});
assign V[86] = {1'b0, V[85][0:126]} ^ (iR & {128{V[85][127]}});
assign V[87] = {1'b0, V[86][0:126]} ^ (iR & {128{V[86][127]}});
assign V[88] = {1'b0, V[87][0:126]} ^ (iR & {128{V[87][127]}});
assign V[89] = {1'b0, V[88][0:126]} ^ (iR & {128{V[88][127]}});
assign V[90] = {1'b0, V[89][0:126]} ^ (iR & {128{V[89][127]}});
assign V[91] = {1'b0, V[90][0:126]} ^ (iR & {128{V[90][127]}});
assign V[92] = {1'b0, V[91][0:126]} ^ (iR & {128{V[91][127]}});
assign V[93] = {1'b0, V[92][0:126]} ^ (iR & {128{V[92][127]}});
assign V[94] = {1'b0, V[93][0:126]} ^ (iR & {128{V[93][127]}});
assign V[95] = {1'b0, V[94][0:126]} ^ (iR & {128{V[94][127]}});
assign V[96] = {1'b0, V[95][0:126]} ^ (iR & {128{V[95][127]}});
assign V[97] = {1'b0, V[96][0:126]} ^ (iR & {128{V[96][127]}});
assign V[98] = {1'b0, V[97][0:126]} ^ (iR & {128{V[97][127]}});
assign V[99] = {1'b0, V[98][0:126]} ^ (iR & {128{V[98][127]}});
assign V[100] = {1'b0, V[99][0:126]} ^ (iR & {128{V[99][127]}});
assign V[101] = {1'b0, V[100][0:126]} ^ (iR & {128{V[100][127]}});
assign V[102] = {1'b0, V[101][0:126]} ^ (iR & {128{V[101][127]}});
assign V[103] = {1'b0, V[102][0:126]} ^ (iR & {128{V[102][127]}});
assign V[104] = {1'b0, V[103][0:126]} ^ (iR & {128{V[103][127]}});
assign V[105] = {1'b0, V[104][0:126]} ^ (iR & {128{V[104][127]}});
assign V[106] = {1'b0, V[105][0:126]} ^ (iR & {128{V[105][127]}});
assign V[107] = {1'b0, V[106][0:126]} ^ (iR & {128{V[106][127]}});
assign V[108] = {1'b0, V[107][0:126]} ^ (iR & {128{V[107][127]}});
assign V[109] = {1'b0, V[108][0:126]} ^ (iR & {128{V[108][127]}});
assign V[110] = {1'b0, V[109][0:126]} ^ (iR & {128{V[109][127]}});
assign V[111] = {1'b0, V[110][0:126]} ^ (iR & {128{V[110][127]}});
assign V[112] = {1'b0, V[111][0:126]} ^ (iR & {128{V[111][127]}});
assign V[113] = {1'b0, V[112][0:126]} ^ (iR & {128{V[112][127]}});
assign V[114] = {1'b0, V[113][0:126]} ^ (iR & {128{V[113][127]}});
assign V[115] = {1'b0, V[114][0:126]} ^ (iR & {128{V[114][127]}});
assign V[116] = {1'b0, V[115][0:126]} ^ (iR & {128{V[115][127]}});
assign V[117] = {1'b0, V[116][0:126]} ^ (iR & {128{V[116][127]}});
assign V[118] = {1'b0, V[117][0:126]} ^ (iR & {128{V[117][127]}});
assign V[119] = {1'b0, V[118][0:126]} ^ (iR & {128{V[118][127]}});
assign V[120] = {1'b0, V[119][0:126]} ^ (iR & {128{V[119][127]}});
assign V[121] = {1'b0, V[120][0:126]} ^ (iR & {128{V[120][127]}});
assign V[122] = {1'b0, V[121][0:126]} ^ (iR & {128{V[121][127]}});
assign V[123] = {1'b0, V[122][0:126]} ^ (iR & {128{V[122][127]}});
assign V[124] = {1'b0, V[123][0:126]} ^ (iR & {128{V[123][127]}});
assign V[125] = {1'b0, V[124][0:126]} ^ (iR & {128{V[124][127]}});
assign V[126] = {1'b0, V[125][0:126]} ^ (iR & {128{V[125][127]}});
assign V[127] = {1'b0, V[126][0:126]} ^ (iR & {128{V[126][127]}});


//assign Z[0] = 128'd0 ^ (V[0] & iCtext[0]);
assign Z[1] =  128'd0 ^ (V[0] & {128{iCtext[0]}});
assign Z[2] = Z[1] ^ (V[1] & {128{iCtext[1]}});
assign Z[3] = Z[2] ^ (V[2] & {128{iCtext[2]}});
assign Z[4] = Z[3] ^ (V[3] & {128{iCtext[3]}});
assign Z[5] = Z[4] ^ (V[4] & {128{iCtext[4]}});
assign Z[6] = Z[5] ^ (V[5] & {128{iCtext[5]}});
assign Z[7] = Z[6] ^ (V[6] & {128{iCtext[6]}});
assign Z[8] = Z[7] ^ (V[7] & {128{iCtext[7]}});
assign Z[9] = Z[8] ^ (V[8] & {128{iCtext[8]}});
assign Z[10] = Z[9] ^ (V[9] & {128{iCtext[9]}});
assign Z[11] = Z[10] ^ (V[10] & {128{iCtext[10]}});
assign Z[12] = Z[11] ^ (V[11] & {128{iCtext[11]}});
assign Z[13] = Z[12] ^ (V[12] & {128{iCtext[12]}});
assign Z[14] = Z[13] ^ (V[13] & {128{iCtext[13]}});
assign Z[15] = Z[14] ^ (V[14] & {128{iCtext[14]}});
assign Z[16] = Z[15] ^ (V[15] & {128{iCtext[15]}});
assign Z[17] = Z[16] ^ (V[16] & {128{iCtext[16]}});
assign Z[18] = Z[17] ^ (V[17] & {128{iCtext[17]}});
assign Z[19] = Z[18] ^ (V[18] & {128{iCtext[18]}});
assign Z[20] = Z[19] ^ (V[19] & {128{iCtext[19]}});
assign Z[21] = Z[20] ^ (V[20] & {128{iCtext[20]}});
assign Z[22] = Z[21] ^ (V[21] & {128{iCtext[21]}});
assign Z[23] = Z[22] ^ (V[22] & {128{iCtext[22]}});
assign Z[24] = Z[23] ^ (V[23] & {128{iCtext[23]}});
assign Z[25] = Z[24] ^ (V[24] & {128{iCtext[24]}});
assign Z[26] = Z[25] ^ (V[25] & {128{iCtext[25]}});
assign Z[27] = Z[26] ^ (V[26] & {128{iCtext[26]}});
assign Z[28] = Z[27] ^ (V[27] & {128{iCtext[27]}});
assign Z[29] = Z[28] ^ (V[28] & {128{iCtext[28]}});
assign Z[30] = Z[29] ^ (V[29] & {128{iCtext[29]}});
assign Z[31] = Z[30] ^ (V[30] & {128{iCtext[30]}});
assign Z[32] = Z[31] ^ (V[31] & {128{iCtext[31]}});
assign Z[33] = Z[32] ^ (V[32] & {128{iCtext[32]}});
assign Z[34] = Z[33] ^ (V[33] & {128{iCtext[33]}});
assign Z[35] = Z[34] ^ (V[34] & {128{iCtext[34]}});
assign Z[36] = Z[35] ^ (V[35] & {128{iCtext[35]}});
assign Z[37] = Z[36] ^ (V[36] & {128{iCtext[36]}});
assign Z[38] = Z[37] ^ (V[37] & {128{iCtext[37]}});
assign Z[39] = Z[38] ^ (V[38] & {128{iCtext[38]}});
assign Z[40] = Z[39] ^ (V[39] & {128{iCtext[39]}});
assign Z[41] = Z[40] ^ (V[40] & {128{iCtext[40]}});
assign Z[42] = Z[41] ^ (V[41] & {128{iCtext[41]}});
assign Z[43] = Z[42] ^ (V[42] & {128{iCtext[42]}});
assign Z[44] = Z[43] ^ (V[43] & {128{iCtext[43]}});
assign Z[45] = Z[44] ^ (V[44] & {128{iCtext[44]}});
assign Z[46] = Z[45] ^ (V[45] & {128{iCtext[45]}});
assign Z[47] = Z[46] ^ (V[46] & {128{iCtext[46]}});
assign Z[48] = Z[47] ^ (V[47] & {128{iCtext[47]}});
assign Z[49] = Z[48] ^ (V[48] & {128{iCtext[48]}});
assign Z[50] = Z[49] ^ (V[49] & {128{iCtext[49]}});
assign Z[51] = Z[50] ^ (V[50] & {128{iCtext[50]}});
assign Z[52] = Z[51] ^ (V[51] & {128{iCtext[51]}});
assign Z[53] = Z[52] ^ (V[52] & {128{iCtext[52]}});
assign Z[54] = Z[53] ^ (V[53] & {128{iCtext[53]}});
assign Z[55] = Z[54] ^ (V[54] & {128{iCtext[54]}});
assign Z[56] = Z[55] ^ (V[55] & {128{iCtext[55]}});
assign Z[57] = Z[56] ^ (V[56] & {128{iCtext[56]}});
assign Z[58] = Z[57] ^ (V[57] & {128{iCtext[57]}});
assign Z[59] = Z[58] ^ (V[58] & {128{iCtext[58]}});
assign Z[60] = Z[59] ^ (V[59] & {128{iCtext[59]}});
assign Z[61] = Z[60] ^ (V[60] & {128{iCtext[60]}});
assign Z[62] = Z[61] ^ (V[61] & {128{iCtext[61]}});
assign Z[63] = Z[62] ^ (V[62] & {128{iCtext[62]}});
assign Z[64] = Z[63] ^ (V[63] & {128{iCtext[63]}});
assign Z[65] = Z[64] ^ (V[64] & {128{iCtext[64]}});
assign Z[66] = Z[65] ^ (V[65] & {128{iCtext[65]}});
assign Z[67] = Z[66] ^ (V[66] & {128{iCtext[66]}});
assign Z[68] = Z[67] ^ (V[67] & {128{iCtext[67]}});
assign Z[69] = Z[68] ^ (V[68] & {128{iCtext[68]}});
assign Z[70] = Z[69] ^ (V[69] & {128{iCtext[69]}});
assign Z[71] = Z[70] ^ (V[70] & {128{iCtext[70]}});
assign Z[72] = Z[71] ^ (V[71] & {128{iCtext[71]}});
assign Z[73] = Z[72] ^ (V[72] & {128{iCtext[72]}});
assign Z[74] = Z[73] ^ (V[73] & {128{iCtext[73]}});
assign Z[75] = Z[74] ^ (V[74] & {128{iCtext[74]}});
assign Z[76] = Z[75] ^ (V[75] & {128{iCtext[75]}});
assign Z[77] = Z[76] ^ (V[76] & {128{iCtext[76]}});
assign Z[78] = Z[77] ^ (V[77] & {128{iCtext[77]}});
assign Z[79] = Z[78] ^ (V[78] & {128{iCtext[78]}});
assign Z[80] = Z[79] ^ (V[79] & {128{iCtext[79]}});
assign Z[81] = Z[80] ^ (V[80] & {128{iCtext[80]}});
assign Z[82] = Z[81] ^ (V[81] & {128{iCtext[81]}});
assign Z[83] = Z[82] ^ (V[82] & {128{iCtext[82]}});
assign Z[84] = Z[83] ^ (V[83] & {128{iCtext[83]}});
assign Z[85] = Z[84] ^ (V[84] & {128{iCtext[84]}});
assign Z[86] = Z[85] ^ (V[85] & {128{iCtext[85]}});
assign Z[87] = Z[86] ^ (V[86] & {128{iCtext[86]}});
assign Z[88] = Z[87] ^ (V[87] & {128{iCtext[87]}});
assign Z[89] = Z[88] ^ (V[88] & {128{iCtext[88]}});
assign Z[90] = Z[89] ^ (V[89] & {128{iCtext[89]}});
assign Z[91] = Z[90] ^ (V[90] & {128{iCtext[90]}});
assign Z[92] = Z[91] ^ (V[91] & {128{iCtext[91]}});
assign Z[93] = Z[92] ^ (V[92] & {128{iCtext[92]}});
assign Z[94] = Z[93] ^ (V[93] & {128{iCtext[93]}});
assign Z[95] = Z[94] ^ (V[94] & {128{iCtext[94]}});
assign Z[96] = Z[95] ^ (V[95] & {128{iCtext[95]}});
assign Z[97] = Z[96] ^ (V[96] & {128{iCtext[96]}});
assign Z[98] = Z[97] ^ (V[97] & {128{iCtext[97]}});
assign Z[99] = Z[98] ^ (V[98] & {128{iCtext[98]}});
assign Z[100] = Z[99] ^ (V[99] & {128{iCtext[99]}});
assign Z[101] = Z[100] ^ (V[100] & {128{iCtext[100]}});
assign Z[102] = Z[101] ^ (V[101] & {128{iCtext[101]}});
assign Z[103] = Z[102] ^ (V[102] & {128{iCtext[102]}});
assign Z[104] = Z[103] ^ (V[103] & {128{iCtext[103]}});
assign Z[105] = Z[104] ^ (V[104] & {128{iCtext[104]}});
assign Z[106] = Z[105] ^ (V[105] & {128{iCtext[105]}});
assign Z[107] = Z[106] ^ (V[106] & {128{iCtext[106]}});
assign Z[108] = Z[107] ^ (V[107] & {128{iCtext[107]}});
assign Z[109] = Z[108] ^ (V[108] & {128{iCtext[108]}});
assign Z[110] = Z[109] ^ (V[109] & {128{iCtext[109]}});
assign Z[111] = Z[110] ^ (V[110] & {128{iCtext[110]}});
assign Z[112] = Z[111] ^ (V[111] & {128{iCtext[111]}});
assign Z[113] = Z[112] ^ (V[112] & {128{iCtext[112]}});
assign Z[114] = Z[113] ^ (V[113] & {128{iCtext[113]}});
assign Z[115] = Z[114] ^ (V[114] & {128{iCtext[114]}});
assign Z[116] = Z[115] ^ (V[115] & {128{iCtext[115]}});
assign Z[117] = Z[116] ^ (V[116] & {128{iCtext[116]}});
assign Z[118] = Z[117] ^ (V[117] & {128{iCtext[117]}});
assign Z[119] = Z[118] ^ (V[118] & {128{iCtext[118]}});
assign Z[120] = Z[119] ^ (V[119] & {128{iCtext[119]}});
assign Z[121] = Z[120] ^ (V[120] & {128{iCtext[120]}});
assign Z[122] = Z[121] ^ (V[121] & {128{iCtext[121]}});
assign Z[123] = Z[122] ^ (V[122] & {128{iCtext[122]}});
assign Z[124] = Z[123] ^ (V[123] & {128{iCtext[123]}});
assign Z[125] = Z[124] ^ (V[124] & {128{iCtext[124]}});
assign Z[126] = Z[125] ^ (V[125] & {128{iCtext[125]}});
assign Z[127] = Z[126] ^ (V[126] & {128{iCtext[126]}});
assign Z[128] = Z[127] ^ (V[127] & {128{iCtext[127]}});

assign oResult = Z[128];

endmodule

