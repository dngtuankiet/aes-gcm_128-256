library verilog;
use verilog.vl_types.all;
entity tb_gfmul is
end tb_gfmul;
